.title KiCad schematic
.include "../models/C2012X7R2A104K125AA_p.mod"
.include "../models/LP38693_ADJ_TRANS.lib"
.include "../models/PCF1C101MCL1GS_v100.lib"
.include "../models/PCF1E100MCL1GS_v100.lib"
XU2 /VIN 0 C2012X7R2A104K125AA_p
XU1 /VIN 0 PCF1E100MCL1GS
R1 /VIN /EN {REN}
V1 /VIN 0 {VSOURCE}
R2 /VOUT /VREF {RADJ}
R3 /VREF 0 {RREF}
XU3 /VIN /VREF /EN /VOUT 0 LP38693_ADJ_TRANS
XU4 /VOUT 0 PCF1C101MCL1GS
I1 /VOUT 0 {ILOAD}
XU5 /VOUT 0 C2012X7R2A104K125AA_p
.end
